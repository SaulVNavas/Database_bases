bit hola
architecture adios
xs if else then fx
aaaa signal
asdfas (library)
www.wait --comments